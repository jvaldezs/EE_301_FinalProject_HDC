--------------------------------------------------------------------------------
-- File: TestHV_RAM.vhd
-- Author: 
-- Date: November 11, 2025
-- Description: 
-- 
-- Revision History:
-- Date          Version     Description
-- 11/11/2025    1.0         Initial creation
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity TestHV_RAM is
    port(
        clk : in STD_LOGIC; -- Clock input from top level clock
        reset : in STD_LOGIC; -- Reset input
        Read_en : in STD_LOGIC; -- Read enable signal FROM THE CONTROLLER/STATE MACHINE
        TestHV_addr : in std_logic_vector(6 downto 0); -- Test Hypervector class address (0-125)
        --controlled by the controller/state machine from bit select module
        bit_addr : in std_logic_vector(7 downto 0); -- Hex digit address (0-255)
        -- controlled by the controller/state machine from bit select module
        data_out : out std_logic_vector(3 downto 0) -- Output 4-bit hex digit
    );
end TestHV_RAM;

architecture Behavioral of TestHV_RAM is

    type RAM_type is array (0 to 127) of std_logic_vector(1023 downto 0);
    signal RAM : RAM_type := (

x"D55C7B6C2DD224E2CBF6286E45715DBC8026AD201B5F36417D577627AC12E6C7C34EBB743248AAEE0E220194BF4EDD96BE861175EA6A7497E9062E905C13DDA0AB074DE5375762E90BFC0303EF5D635F63D1963919713C65C538C3B924884A27B0BCE2C1D9E126131581AF900366485C7340B677E0CD94AA8D5C622094DA95E7", 
x"B54C6F2CADF2A4E38AD6187C4F715F2C8006BD601B5F2161795F36372C92E6E7C34DFB553248ABEE5E2241E6BF4E4D863E871165C063F497ED043C8C4C5B1DA0AB074D85375762E9ABDC4311AF59735973D1D63819717D4FC730C3B864A84E17B01CE2C1C9E1261B1081AF90136EC85473C1B67748CD14A2855866139CDA15E7", 
x"D7CC6F2CAD92A4E34AF6387C07715D3C8016AD219B5F20617D533636AC92A6E7C26BF77132482BEE1EA241C6BE4E4D86BE87517DE262FC97AD062CC85C5FDDA5A32759C53F5622E92BFC4311AF59635973D5963818713D45C53082B86C82C657B09CE2C19DE0261B19032E900376C85473C1F6E758CD14E28578626B9CDA95E3", 
x"C55C4F6E2DF224E3CBF6387C65715D3C8006AD201B5F3541791736222C92E6E7D24EFB513248ABE60F2201C4BF4ECD86BE865575E263FC95A90638D45C1BDDA4AB074DC53F5726E92BFC0311AF59635D63C5D6B809F13D45C330C3B924AACE33B03CE241D9E1261B15812B90136EC8D473C0B667E0CD14A28D5C620BDCDA95E3", 
x"D74C6F6E2DF224E3CBD6286EC5715D1C8032AD60395F3761595776326C1266C7C24FFF503248ABEE0F2240CCBE4E05863E871165E8627497ED063C805C179DA0AB274DA5275E32E98FF04301EB5D635D73D6D63818717D45C138C2B86CA84F03B034E2C1D9E1261B3501AB901366485C7340B27760CD14E28550623394DA95C3", 
x"8BCC4B2C25B224E3CBD638EC07714D3C8022AD205B5F30617F5776372C92A6E7D24AFB503248ABEE1F2241C4AF06CD86BE861165E26BF497ED0408D05C171DA1AB0749C73F5F22E96BFC230BAF5D635D73D1963119713D45C730C3B96C82C633B01C6261D9E1261B3D89AE90137EC8D47140B6E740CD14A28D74624394DA15EB", 
x"B3CC6F3C259224E3CBD6187E47715F3C9026BD601B5F0061595F36066C92E6C7C27AFF503248ABE61F226086BE460D96BE861165E260FC95AD043CC05C1B1DA1A3064DA7234F62E9EBF46301AB5D7359F3D5963918F13D4DC33082B96CA8CE53B01C62C19DE0261331812E801366C87471C1F6F760CD14E28D5C666A9CDA11A3", 
x"915C6F2CADD224E34BD6187C07715D3C8006AD201B5F31615C5776126C92E6E7C24ABF513248AAE61F2240ACAF0E4D96BE861175E26BB497A90420D45C1B5DA1A3265DC7374F63E9AFFC2301AF4D635DE3D5963819713D67C33082BD64A84757B01C624199E1261B1581AE901766C8747342F6E760CD14A2857C627BDCDA95AB", 
x"D75E6F6C85D2A4E38AD6387E85715DAC8006AD619B5F37415B533622EC92E6C7D24DB75032482BEE0F2280A4BF0E05863E865F65E263FC97A9063ED0DC1B5DA0AB264DA5275777E90FFC0301AB59735973D4D63018F13C67C530C2F92CA84733B09EEAC1D9E1261B11012A80037EC8547353B67750CD14A29D58620AD4D21587", 
x"D1CE6F2C2DB2A4E3CBD6187C47714D3C8026BD215B5F04615D5336162C92A667C25ABF513048ABE61F2261A4AF064D96BE86116DE261F495AD063CD05C1F0DA0A30749E7235F2AF92BF82309AF497359F3D1D6390871BC45C33082B064A8CF53B01D62C1BDE126133C812E941376C8747340F6E7E0DD14A2CD74647BDCDA91A3", 
x"F5CE673CADD224E2CBD6386C27615F3C9036AD601B5F11617B5736262C92A6C7C36CB7503248ABE61E2261A6BB4E0D963E86536DE2627497ED0424984C175DA3AB064DE5275F6BE9ABF44301AF59735963D1963909F13D45C730C2B86CA04E57B034E2C1DDE1261318812A900276487C73C0F6F7C0DD14A28D58627BDCDA91A7", 
x"C5DC5F2C2DB224E30BD638FE07F15F2C8006AD60BB5F344179573632EC9266CFD25DF7153048ABEE0E22C0A4BF4E5D863E871165E062B497AD0604C45C1359A6AB074D05377766E92BFC0301AF59735D73C596B819F19D47C138C2F96CAACF52B01CEAC1C9E1261B1901AE90127E48547342F66740CD14A29D5866129CDA15A3", 
x"D5CC6F2CADF224E3CBD6187C67715D3C8036AD211B5F01617F1336162C92A6E7D25ABF513048ABE61F2241A4BE06C596AE86516DE269F495AD043CD05C1F4DA0A30649E53B5F2AE92BF86309AF4D6359E3D1D63918713D47D738C2F92CA2CF53B01C62E199E126131C832F941376C8F47140F6E7F8DD14EA8D5C647BDCDA11A7", 
x"D55E6F2CADF2A4E34AD6387C05715D3C8002AD201B5F23617D5736172C92A6E7C24FF7553048ABEE0F2240E4AF0E5D86BE86516DE2637497E9063CD85C575DA4AB075DE53F5662E92FFC630BAF4D635D73D5963818F13D45D73082B92488C637B09C62C19DE0261315012F90137E485471C0B6E7D0CD14E28D58727BDCDA95EB", 
x"D54C6F2CADF2A4E3CBF6386C67715F3C8002AD601B5F354179577626AC92A6C7D25EB7543248ABEE1F2240C4BB4ECD963E87517DE26BF497ED063CC84C179DA0AB024DC53B4E66E9ABFC4301EF59735F73D5D63818F13C4DD338C3B92C88CE15B01CE2C1D9E126131581AF900376C87C7341B6E740CD14A28D78620ADCDA95E3", 
x"D55C4F2DADD2A4E3CBD638FC45715D0C8016AD611B7F374179533603EC92E2E7D37FB7313248ABE64E22E1CEBF4E05863E871165E263BCB5E9041ED4DC1F9DA0AB064DA5377E27E9EBF8030BAF59735B73D5963009713D45C730C2B924AA4F13B09C62C1D9E1261311032F90027EC85C7352B66760CD14E29D787262D4DA15E3", 
x"C54E5F6E2DB2A4E3CAD6386E47715D2C8026AD20FB5F014179173633EC92E2E7D36CBF3032482BEE0F2201A4AB0E1D96BE865965F06BF4B7A9041CD4DC179DA1A3074D873F5F27E9ABF82309AF59635B63C5963818717D45C73083B96C80C631B01CE2C1F9E1261B1903AD90036EC85C7340F6E740CD14E285786243DCDA1583", 
x"955C6F2CADD224E3CBD6286C05715D3C8032AD603B5F2561791736026C92A2C7D24EBB713248AAEE0F2240D4BE4EC586BE871365E2637495ED062ED05C575DA0AB274DC5275F32E9EBDC230BEF5973DD73D7D43818713C45C138C2B964AACF13B01462C199E1261B1D01AA801376487C7340F66760CD14A28D50625A94DA95E3", 
x"85DC6F3CADD224E3CBD6186E67715D3C8026AD21F95F214159573602AC9266E7D25EB7503248ABEE0FA241C6BE4E0D96BE865165E262BC95ED063C904C1F99A0AB034DE76F5F72E90BD86301AB59735BE351D43908717D47C13882B96C88C671B03F6241FDE126173C812F901766485C7340B6E7E8CD14AA8D74642BDCDA91E3", 
x"F5CE4F6CA5B2A4E3CBD6186C67715D3C8026BD203B5F2161795F36162C92A647D258BF513248ABEE1F22C0A6BA4E0D96BE861165F260FC95AD043CD8DC1F4DA0AB0749876F5F76F90BF02303AF4D735963D7D43908713D47C330C3B82CA8CF33B01C62619DE126131C81AE801766C87473C0F6E7685D14A28D78644A9CDA91E7", 
x"854C6F2D2DF224E34BD6386C67715D3C8036AD207B5F31615F5776366C92A6E7C34AFF513248ABEE4F2241CEBB4ECD863E86517DE261F495ED062CD05C1FD9A1A30659C5335E76E96BF86301EF49735973D5963819713C45C730C2B82CAACA73B015E2C1D9E1261B1001AE901366C8747141B6E740CD14EA8578722BD4DA15C3", 
x"95CC4B6D2DB2A4E30AD6386C67715F3C8012AD201B5F31617F573632AC92E6C7C24AFF513248ABEE1FA241E6BB4E4D86BE861175C263F497ED060CD85C171DA5AB275DC5375F27E92BFC4301EF59735B734196B819F13D67C730C2B96C824673B01FE2C1D9E0261B1C032A90136EC85473C0B677C0CD14E28D78606B9CDA118B", 
x"D55C6F2EADF224E3CBD6286C25615D8C8012AD205B5F25417B177636AC9226C7D24FFF503248AAEE0E2260C4BF0EC5863E87116DE263F497ED062ED04C175DA5AB074DC5376776E9CBDC0301EF59635D73D5D63819713D65C738C3B924AACE37B01462E1D9E1261B15012E901366C85C7300B66670CD14A28D50626A94DA15E3", 
x"D5DC6F2CADD224E34BD6386E05715D3C8022AD201B5F204179577636AC92E6C7D34AFF513248AAEE0E224084BF4EC586BE061365E263F497ED062C90DC1F1DA0AB074DC5374E76E90BF84301AF59635DF3D5D63819717C45C738C2B92CAA4E15B01C6241F9E1261B11012E901366C87C7340B6E768CD14A28D50666BD4DA95E3", 
x"855E4B3CAD92A4E34BF6386C67715D3C8012AD201B5F20617B533626AC92A6E7C24AFF503048ABEE0F2241C4BF06C596BE86116DE22BBC97E90634905C139DA0A3064DE5275F7FE98BF84301AF59735973D5963919713C45C73082B96C88CE13B01CE241DDE126131581AE801366C87C7340B6F760CD14AA8D58626BD4DA95E3", 
x"975C5B2EADD224E34BD6286C07F14D2C8006AD60BB5F3761591776232C92E6CFD24FF3543248ABEE1E224094AF0E4586FE87557DE2617495E9022E945C1FDDA0AB0749E5277F67E90BF82303EF5D635B73D5963119713C45C730C2B924884F17B094E241D9E1261B1509AF840366405C71C0F26760CD14A29D54667A9CDA95E3", 
x"D54C4F2C25D2A4E2CBD6387C47715F1C9026AD603B5F0141791F3636EC9266E7C26BB3513048ABEE1F2240C4AF4E4D963E86516DE260FC97ED0438C85C175DA1A3074987335B23E92BF44303EF49635963D5D63919F19D4DC730C3B82482CE73B01C62C1F9E1261B1501AA90127E485471C0B2E770CD14E28574665ADCDA95E3", 
x"D55C7F2C25F224E3CAD6286C67715D0C8006AD203B5B37617A1736322C1266C7D34FFF7532482BEE4E2240C4BF4E0D86AE875565E063F497E9043CD05C1F9DA4AB0749E73F6777E9EBF8030BAF5D735F63D5D63909F17D45C538C3B92CA84F13B01CE241DDE1261B11812F80136EC05C73C0F67778CD14A28D5C6618DCDA15E3", 
x"854C6B2E2DD224E24BD6387C67615F1C9016AD603B5F01617F5F36222C92E6E7D278F7703048ABEE1FA241EEBF4E45963E861165C2637C97E9043C984C1F8DA5A32259853F7726E90BF44309AF59635973D5D63818713D4FC53083BC6CA2C633B03DE2C1D9E0261310012E90027E485C7380F6F6C8ED14E28D54646A9CDA95EB", 
x"D74E4B6EA592A4E2CAD6387E47715D3C8006AD201B5F0041585736062C92A647C358F3113248ABEE0F2241C4BE4ECD96BE865365E229FC95ED043C944C5F0DA1A3024DC5235726E92BFC230BAF49335BE355963818713C47C13082B96C884753B01C62E1D9E126171401AE80167EC87471C0F6F760CD14A2CD7C646A9CDA91A3", 
x"C74C6F6C2DF224E34AF638FC05715D2C9026AD20195F34417C5776276C92E6C7C24FBF513248ABEE0E2240DCAE0E1D96BE861165CA62F497E9042CCC5C175DA1AB274DC5374F37E98BF84309AF4D635973D1963819F1BD45C530C2B92CA24773B09CE2C1D9E0261B19012E90027EC85473C1F6E7C0CD14A28570624BDCDA15A3", 
x"D5CC6F6C25D224E2C3D6386C47715F3C9026BD203B5B04617D573626AC92A6E7C35AB3503048ABEE4F2241AEBA464D96BE861175E061FC97AD0638D84C171DA1A30649C7275F6AE92BF82313AF5D3359E3D1D43908F13D45C738C3BC6C8ACF13B01C62C199E1261B3401AE80177EC87471C1F6E740DD14E28D74644BDCDA11AB", 
x"87CC7B2C25F224E3CBD6286EC5714D2C8006AD20795F37617D577617AC9266C7C34AF75532482BE64F22C0E4BF4ECD86BE861165C0627C95E9063CC4DC1B59A0AB264D053F5E76E96BF80301AF5D735D6351D6B919713C67C53882B96CAA4E15B01CEAC1B9E1261B1D832B941366405473C0F66770CD14A28D5C7A1BD4DA95E3", 
x"C74C6F7CADF224E3CBD6386C25715F1C8006BD203B5F21615F5736162C1226C7C24EFF503248ABEE4F2240CCBA4E4D863E875165CA69F497ED063CC05C1F5DA5AB065985377F36E92BFC4301EF5933597351D63908713D45C53082BC2CAACE73B01C62C1DDE1261B1901AF901376C8547140B6E7F8DD14EA8D786203DCDA15E7", 
x"D5CC6F2C2DD2A4E24AD6186C47715D3C8006AD605B5F21617D573626EC92A6E7C25BB7503048ABEE5F2241C4BB4E0D96BE861165E223F497ED063C9C4C174DA1A3024DE7635E66E94BFC630BAF5D335DF3D5943119717C47C530C3B16CA84743B01462E1D9E1261B35012E80177EC8747181F6E7C0DD14A2CD58606BDCDA11E3", 
x"85DC472E2DD224E3CBD6286C45F15D2C8022AD60795F356178577622AC92E6C7C24EB3553248ABEE0E2240A4BF4E0D86AE86137DEA63F497A9043ED45C175DA2AB0749273F6767E9CBF0030BAF5D635DF355D63009F13C67D130C2B924A04F37B09CE2C1D9E1261B1181AE800776485C7340B6F7E0CD14A28D547233DCDA95E3", 
x"87CC6F6D2DD224E3CBD6287EC7F15D0C8012AD601B5F27617A1F7633AC1266E7C34EBF5030482BEE0F2201A4BF4E9D863E87116DE063F495E9060CC45C179DA1AB264D85375777E92FF80309EF5D73597355D6B819711D67D538C2B82C824E21B09CE2C1F9E1261B1581AF901366405C7380B66770CD14E28D58760294DA95E3", 
x"875C6F2C2DB2A4E34AD6386C25715D3C8006AD201B5F3141795776332C92E6E7C24AFF5132482BEE0F2261E4BF0EC586BE865165E262F497ED043CD05C171DA7AB0659E53F5F36E90BF84303EF5D635973D1963008713C45C538C2B82CA24653B01D6AC1D9E1261B1901AA90137EC8D47342B6F758DD14AACD58626ADCDA11E3", 
x"D75C6B6EADD224E3CBF6186C25715D3C8026AD211B5F364179177622AC92E6E7D24FFF753248ABEE0F2241D4BF4E0596BE861775E26AF495E90620D45C139DA0AB074DE53F567EE98BF86303AF5D63DD73D5D63019713D65D530C3B924A2CF07B03C6241D9E1261B15812E800366485C7340B67770CD14A28D5C622394DA95E3", 
x"C55C5F6CA59224E24BD6286C07715D2C8022AD605B5F2561781776222C1266C7D34BF3503248ABEE4F2200C4AF0E4D96BE87157DE26BF495ED0622D45C17CDA0AB074DE5375637E90BF8230BEF5D635B73D7963119713C45C330C3B86CAACF23B01CE2C1D9E1261B1581AF801766485C7340F677E0CD14A28D7C607B94DA15A3", 
x"D14C6B6CADF224E34BD6186C07715D3C8004AD601B5F04617F5336062C92A6E7D24ABF513248ABE64F220184AA464596EE865165E2687C95ED063C904C1B09A1A3034DC5275F3EE90BFC0311AF4D3359E351963119F13D45C13083BD6CA24F43B01C62C1FDE1261310012E90167EC85C7140F6F760CD14AADD706469DCDA91A3", 
x"95CC6F2D2DB224E2CBD6286EC7715D2C8022AD603B5F25617B5B3636AC92E6C7C34FF71030482AE64EA24084AE0E4D86BE865165C2607497ED0624C85C534DA5AB274D85375E26E92BDC4301EF59635973D7963019713D47C53883BC6C8AC665B09CEAE1D9E1261B1401AE901376485473C2B66748CD14E2857876139CDA91E3", 
x"97DC6F6CADD2A4E3CBF6287E45715D3C8016AD201B5F356179577623EC92E6C7C25EFB553248ABE64F224184BF4EC596BE861165E262F495E90634D05C179DA0AB074D65275626E98BF84303AF5D635D73D1963818717D45C738C3B964A2CE13B09C6241D9E1261B11012B900366487C7340B667F0CD14E28D50667B9CDA95E3", 
x"87DC7F6E25F2A4E3CAD638FE67715D1C8026AD60395F3141791F36336C9AE2E7D34FFF3032482BEE0E2200E4BB4E0D963E865565EA6BB495E90408DCCC175DA7AB274DC5274766E92FF82301EF5963D963C5963908717D4FC730C3B92C82C213B01C6AE1D9E0261B3101AD90136E485473C3B6E7D0ED14A2857C60429CDA15C3", 
x"D55C6F6EADF2A4E3CBF6287E67715D0C8002AD411B5F37417B1736132C92E6E7D35EFB743248ABEE0F220184BF4E8D963E87196DEA63FC97ED062E984C170DA2AB074D85377667E9CBD80311EF59735963D5963108F17D65C730C2B824AACE23B0BC6AC1D9E1261B11012F90136648547341B67768CD14E28D58626B9CDA95E7", 
x"D14E6B2DADF2A4E3CBD6187C27715D3C8012AD201B5F24615F5736062C92A6E7C25AB7513248ABE61F224084BB060D96AE865965E269F495ED063CD05C1F1DA1A32349E5335F2EF90BF4630BAF497359E3D5D63918713C47D33083BD6CA8CF13B01D62419DE1261319812E80176EC8F47340F6E768DD14EADD7C647B9CDA11A3", 
x"954E6F6E2DF2A4E3CBD6386E25715D1C8032BD611B5F31617F5F36362C1226E7C24BF7113248ABEE4F2240C4AE4E4D863E861165E261FC97ED0430C85C17DDA5AB065DA5375E26E92BF86303AF5D73597351963008717C45C530C3BC6C884E73B01C6241DDE126131101AA901376C8547180B667C0DD14AA8D78600B9CDA15E3", 
x"874C6F3CADB224E3CAD6386C67715D3C9002AD211B5F31617D5F76372C9226C7C24EF75132482BEE0F2260E6BF4E4D86BE871165E269B497ED0604C05C17DDA0AB025D85375F76E90BFC6301EF59635973D596B918F15C47D738C2F92CA8CE13B01DE241DDE1261B1981AE90136EC85471C2B6E7C0DD14EA8D78622BDCDA15A3", 
x"D7CE6F2CA592A4E3CBD6187E07711D3C8006AD21795F34617B5776372C9222E7C24AFF5032482BEE0FA240A4BB464D962E865965E26AB495ED0428C05C135DA1AB274DE53F4F66E96FF04301AF59635963D596391871BD47C33083BC6CA8CE53B01C62419DE026131581AF901366C8547142B6E760CD14AACD746E6B9CDA95A3", 
x"C54C5F2D2DF2A4E3CBF6386E47F15D2C9026AD201B5F34617C5336332C92E6C7C34FFF113048AAEE0F2241A4BF4E0D863E861565E022F495E9062CCCDC175DA7AB275D45335E66E92FFC0301ED5D735D7355963018F15D47C530C2F86C0AC631B01C62C1D9E0261B3981AE900366C8D473C2B67740CD14A29578721394DA15C3", 
x"D5CC6B6EADD224E34BD6386E45715D0C9012AD60BB5F356179173637AC92E6C7D34FFF7132482BEE4E2281C4AE4ECD863E86116DE26B7497E9063EC45C1F1DA6AB064D8537763FF90BD04301AB59735D73D5963019F13C45D530C2BC6CA0CE07B01CEAC1DDE1261B1D01AF90136E405C7350B67760DD14E29D5C620BD4DA95E3", 
x"F1CC6B2CADF2A4E24AD6187C67710D3C9026AD203B5F24615F5336062C92E6E7C24AB7503248ABEE1F2241A6BF460D96BE861175E268FC95A9043CD45C1F1DA1A32649C53B4F22E9ABF42309AB5D335973D1963919713D67D33082B96CAA4F57B01D626199E026131181AA901676C87471C3B6E7E8CD14A2DD7064639CDA91A3", 
x"D5CC6F3C2DF2A4E3CAD6386E47715D3C8022AD20BB5F31617B5376262C9226E7C24AF3503248ABEE4F2240A4AF0E4D86BE86517DE263F497AD042CD45C1BDDA0AB0749C73F4E22E90BF04303AF4D635B73D5963818713C47D738C3BD2482C613B01CE2C19DE1261B3581AE901366C85473C0B6E7E8DD14A28D5462739CDA95E7", 
x"D55C6F7DADF224E3C3D628EC47715D1C8022AD21795F3561795776326C1266C7C34EFF5032482AEE4FA260C4BF4ECD86BE871165C862FCB5ED0420C05C174DA0AB274D853F6E6FE9AFF82311EF5D635D73D796301871BC47D330C3B864AACE07B03462C199E1261B1981AF901366485C7150B66768CD14A28570625B94DA1583", 
x"F34C6F2CA5F224E3CAD6187C25715D3C8026BD20195F30615F5736062C92A6E7D24ABF503248ABEE0E2261A4BB464D96BE86116DF263F497AD063CD05C1B19A0A32649E7335F66E9EBFC6309AF5D735BF3D1963918F13D65D730C2BD2CAA4753B09C62C19DE0261311012E901376C85473C2F6E7E0CD14A2855C6463DCDA11A3", 
x"F7CC6F2CADF224E3CBD6187C67715D3C8006AD217B5F2161795B76062C92A6E7C25ABF513248ABEE4F2241A6AF0E4D96BE865175E268F497AD043CC05C1B4DA1AB0749C7375F22E92FF82313AB4D735BE3D1D63918713D47D530C2B86C8ACF73B01D62E19DE126131181AE901776C8D471C0B6F7E8DD14AA9D7C647ADCDA95A3", 
x"9D5C6F2DADB2A4E3CAD6387E45715D3C8022AD205B5F2041795376326C92E6E7C26FB71532482BEE0F2241B4BE4E4D86BE861165E2637CB7E9042CC45C1359A6AB074DA5377276E9EBF04309EF5D635F73D596B818F13D45C538C2B824A04753B01EE241D9E1261B19012E90137EC8DC73C0B66740DD14E28D5C6242DCDA15A3", 
x"87CC4F3DADF224E38BD6386E47715D3C9002AD61B95F35415D5736166C9266C7C35EFF1132482BE60F2280F4BB0E4D963E87196DEA603C95ED0638C0DC5F9DA3AB264D85375E6FE92FF80309AF5D735DF3D7963809793D47D53882B86CAA4E07B0B4E2419DE1261B3D03AE90136EC8547140B66640CD14E29574721A94DA95C3", 
x"D94C4F2EADF2A4E34BD6086C65F15D2C8032AD211B5F31415D1376062C9266E7C25AFF503248ABE60F2251ECBA46C586BE86116DEA6AFC95ED041CD04C1F0DA1AB264DC5275E77E9CBFC6301AF59635DE3D1D63908713C47D33882B96CA8CE13B0146261D9E126131581AE901366C87C7102B677604D14E28D5C626394DA15EB", 
x"C5DE6F3CADD2A4E3CBD6386CE7715D1C8012AD201B5F31615B5736332C92E6C7C34AF7503248ABEE1FA200C4BF4E4D863E865167E260FC97AD0634D45C175DA7AB264D853F576EE94BF06303AF5D735973D596B118713C47C738C2B96C8A4E31B03462C1D9E1261B1501AE90137EC87471C0B6E7C0DD14EA8D7862339CDA1583", 
x"D5CC7B6CADD224E3CBD6286E05715D2C8006AD00FB5F34417D177632AC1266C7C34FFF1132482BEE0E22C1C4BF0E4D86BE861165EA62FC97E9042CCCDC1F5DA0AB065DE5377627E9ABF40301EF59235F73D5D63919715C45C538C2FD6CA84703B09CE241D9E1261B1981AF90136640547342B66760CD14EA8D586E1294DA95A3", 
x"855C6B6CA5F2A4E3CBD6387E47715D0C9002AD60997F3141595776336C12E6E7D24EBF113248ABEE4F2201E4BF4E4D863E871165E261BC97E90628C4DC575DA1AB064D85377F77E9CBFC030BEF5D735D73D5963808F17D45C730C2B824AA4E23B01CE2C1D9E126131101AE900366C0547342B6F740DD14E29558720894DA15E3", 
x"95CE6F2CADB2A4E3CBD6186C67715F3C8026BD203B5F30617B1736166C92A6E7C24ABF113248ABE61FA241ECBA460D96AE861165E261B497AD043CD0DC5B4DA1AB024DC7335F26F96BFC2309AF59735D73D596391871BD45C13082FC2CAACE13B03C6261B9E126133501AE901376C8DC71C1B6F7F0CD14A2DD7C6469DCDA11A7", 
x"955E6B2C2DD224E34BD6286C65715D1C8002AD201B5F224178537633AC92E6C7D34EFF303248AAEE0FA240E4BF4EC586AE87516DE2607495E9043CD05C575DA0AB034D85375677E90BD80311EF5D23DD73D4963108793C47C738C3B964824E17B094E2C1D9E1261B1D01AE90136648547342B667C8DD14E28558722B94DA15C7", 
x"D55C6F6EAD9224E3CBF6386C65715DBC8016AD601B5F31617A5F76126C9226C7D34EFF553248ABE60E220084BF4ECD867E871165E26BFC97E9062EC05C131DA1AB075DC5377736E90BFC0303EF59735F73D5D63009793D45C53883B824A84E37B09C6241D9E1261B1181AF901376C85C7340B67778CD14A28D58623B94DA95E3", 
x"D5CC6F2CA592A4E24BD6186C27715F3C8016AD201B5F00615F1776162C92A6C7C26AFF113048ABE60F2241A4AE06CD96BE865165E269F497AD042C905C171DA1A30749E5375F22E9ABF46309AF5D3359F3D196381971BC45C330C2B86488CF33B01F62419DE126131181AE90176EC8F47140F6F760DD14E29D74647ADCDA11A3", 
x"C55C7B2CADF224E3CBD6286C27715D2C9002AD20F95F30617B5776322C92A6E7D34EFB513248ABEE0F224184BF4E8D86BE861575EA6BBC95ED062AD45C13DDA5AB074DE73B4F66E94BF0031BAF5D235B73D596B009F13C47C730C3B964A24F63B01C62C1D9E1261B1D81AF90136648D473C0B66768CD14A28D7862589CDA15E3", 
x"C55E433DAD9224E2C3D6386C67715D3C8036AD603B5B21617B573636EC92E6E7C359F3503048AAEE1FA240CEBE4E4D96BE865365E223FC97ED043C984C1F0DA1A3274DC72F4F2EE92BFC630BAF5D735BF351963119713C47C138C3B96CAA4753B0956241D9E0261F1D81AA94127648747300F6E740CD14E2CD5C645A9CDA11EB", 
x"D55C4F6C2DF2A4E3CAD6286C47715D2C8016BD219B5F2341795736332C92E6E7D34FF75532482BEE0F2220C4BF4E1D863E861165E262F4B5ED042CD05C17DDA0AB2749873F5F66E96BF80309AF5D735D73D1D6B019F17C45D730C2B82CAAC613B01E6241D9E1261B15812F90037EC8747140B667E0CD14E28D70625B9CDA11A3", 
x"95CE4B3CADF224E2CBD6186C27715D3C8026BD205B5F20617F1336162C92A6E7C26AFF513248ABE61F224184B7464D963E86116DE229BC97A90638D0DC571DA1A3064DC5335F6FF98BFC631BAF597359E3D1963818713D47C530C2B92CAA4E13B01E6261DDE126131D012E80137EC8D471C1B6E7E0CD14E29D5C6462DCDA15E3", 
x"C54C477CADB2A4E3CBF6387C47715D3C8026BD201B5F21617B573626AC92E6E7C24AF3503248ABEE1F2241A4BF4E4D96BE865175E263F497ED042CD85C1F1DA1A30649A5375F72E9EBFC6311AF59735963D1943818F13D47D738C2B96CAAC673B01C62C19DE1261310012F90137EC85473C1BEF7E0CD14E28D746263DCDA11E3", 
x"DD4C672CAD92A4E2CBD6186C67615F3C9014AD213B5F31417B573622AC92E6E7C36CB7503248ABEE0F2251A6BB0E4D963E865165C26BF497ED0434885C175DA1AB064DE7236F3EE9CBFC2311AF493359F351963918713C45C538C2B96482C657B0BDEAC1DDE1261310012A900676487473C1F6F7C0CD14A28D74626ADCDA91A7", 
x"D55C4B2CADF2A4E34AD6287C45715D2C8026AD20BB5F23417D573632AC9266C7D35EFB553248ABEE0E2260F4AF4E4D863E86156DEA63F495E9043480DC135DA2AB064DE5334F67E94BFC030BAF59635963D1963819F13C45D530C3B82C80CE17B01CE2C199E1261319012E901376487473C0B67760CD14E29D5C6212DCDA15E3", 
x"85CC6F2C25F2A4E24BD6187C07715D3C9026AD20BB5F05417B573602AC9226E7C24CFB553248ABEE1F2260A4BF0E0D863E865565E263F495E90424C05C131DA0A32759C7337E67E92BF80309AF5D735973D1943819F13D47C530C2B864A8C217B01CE2C19DE1261334812E801276C85471C0B6E740DD14AA857462729CDA95A3", 
x"855C6F3E2DD224E3CBD6286EC5715D0C8022AD203B5F2741795F7633EC12E6C7C34FFF1132482AEE4F2240ECBE4E45863E87116DC062F4B7ED06288CDC1F9DA2AB274DA737466EE98BD8030BEB5D635D63D7D6B919717D47C138C2B864AACE17B0946AC1B9E1261B35012F901766487C7340B66760CD14E28550663B94DA95E3", 
x"C75C6F2CADD224E3CBD6386E25715DAC9026AD201B5F3461595736062C92E6E7D24FF3343248ABE61E2261DCAF0E4D86BE86116DC22BB497E90628DC5C1F5DA3AB0649E537563FE9ABFC6309EF59635B7351963818713D45C730C3B964A04E17B01CE2C1D9E1261311012F90136E405C7342B67740CD14A28D586243DCDA95E3", 
x"95CE6F2C2DD2A4E3CBD6386E65715D2C8412AD60BB5F25415B577637AC1266C7D25BFF1032482AE60E2200CCAF4EC5863E86116DE263F497ED063CC8DC17D9A7AB235DC5335E7FE98FFC4303EB5D735D73D596B818797C55D738C2B82C8ACE03B0BCE261CDE1261F1983AF901366C85C73C0B66740CD14E29558622B94DA95CB", 
x"D54C4B2C2DD224E34BD6386E07715D3C8022AD61195F004179173636EC9AA6E7C34FB71132482AEE0F2281A4AB4E0D96BE871175E263F497E9063CD44C530DA0AB064DC53F562EE9ABF84309AF59635F63D5D63819F13D45D538C3B82CAA4E03B01C62E1D9E1261B11012F90137EC07473C0B66740CD14E28D70761ADCDA15E3", 
x"955C6F7EAD9224E2CBD6186C47715D3C8006AD201B5F206179573612AC92A667C34AFB553048ABE60FA240A4BE464D96AE865575C263FC95ED063CD04C170DA1A3264DE72B4F26E96BF86303AF59335BE351963119713C45C7B083BC6CA0C643B0146241D9E126133D012F90167EC8547140F6F7E0DD14A29D5C64709CDA95A3", 
x"D54C6F2DADF2A4E38AD6387E45715D2C9022AD613B5F11417F5776336C9266E7D24FFF143248ABEE0F2260C4AF0E1D863E86516DC261FC95ED062CC45C1B5DA1AB274DC5235E66E92BD06303EF5D735973D5D63819F1BD4FC730C2B86CA0C713B03DE24199E1261311832F900366C85C73C0F66748CD14E2C578620A9CDA15A3", 
x"915C6F2E2DD2A4E34BD6287CA5715D2C8006AD609B5F31417D5736336C9266E7D24FBF103248ABEE0F2240C4AF0E1D863E87516DCA62F497E9062ED84C1FDDA4AB275985337627E94FDC4303AF59635973D5D63818717C4DC730C2BD24A2C637B09E6AC1D9E126131503AF90136648547302B67760DD94A28558624B9CDA15C3", 
x"C15C6F3C2DF2A4E2CAD6386C47714D3C8006AD21F95B2461795736322C92A6E7C258B7503048ABEE4F2241ECAA461D96BE865575F262F497E9043CD84C174DA1AB0349C76B5F2EE92BF0630BAF4D335B73C3D43919717D47C53083BD6C82CF13B015E241D9E126171501AE801276C8747140F6F7E0CD14A28D7C746ADCDA95A3", 
x"D75E6B6CADB224E3CBD6386C25715D1C8022AD203B5F34417D5736122C1226E7D25ABF553248ABEE4F2240CCBF4E45863E86536DE223FC95E9063CD04C1F9DA5AB034DC52F5F32E9ABFC2303EF59735F73D5D6381871BC45C338C2B96C82CE13B03D6241D9E1261B1501AF901376C8547140B2F750CD14AA8D5C666B9CDA15E3", 
x"95CC7F2CADF224E34BD6386E45715D2C9022AD603B5F35417F533637AC9266C7C24BFF5132482BEE0F2280E4AF4E0D963E87156DC862FC95ED062CCC5C1759A1AB275D85377F67E96BF80301AB5D7359F3D596301879BD47C130C2B96C8AC633B01CEAC19DE0261B1001AE90036EC8547380B6F740CD14E28D5C761B9CDA1583", 
x"D5DC4F2CADD224E3CBD6386C65715D3C8002AD201B5F31417B5776322C92A6C7C34EF75032482BEE0E2201C4BF4EC5863E86517DE2637C97E90624D45C575DA0AB274DC53B5F27E9CFD80303EF5D635973D5963818713D45C730C2B96488CE17B01EE2C1FDE1261B19812B901376C85C7140B667D0CD14A28558626B94DA15E3", 
x"99CE6F2CADD224E24BD6186C47715D1C8016BD201B5F30615F1376162C92E6C7C25AFF513248ABEE0F2261C4AE064D96FE86516DE269B495AD043CD45C535DA2A30649E7375F2AE9EBF82301AF4D7359F3D5963818713D4DD338C2B92CAACF73B01D624199E1261319012E841766C8F47100F6E768DD14A28D7C667ADCDA15A7", 
x"934C6F3CA5F2A4E2CBD638FE65715F1C8006BD601B5F21617B5736262C92A6E7D37EBF503048ABEE5F2241F6BF0E4D963E86136DE262F497E90434885C1F9DA0A3074D87776726E92BFC430BEF5963596355963819F17D4DC53882B864A2C733B014E2C1D9E126171181AE801276C85473C1F2E7C8CD14E28574622A9CDA95AB", 
x"D55C6F2D2DB224E3CBD6386E45615D3C8022AD013B5F24417B537633EC1226C7C34BBF5132482AEE0F2241C4BF4E45863E875175E2627C97ED0424D05C535DA0AB275DC5377F36E94BF82303EF59635F73D1963008713C45C738C3B924A8CE05B01662C1D9E1261B1D812E900366C85C7340B6E740CD14E28558626BD4DA15A3", 
x"975C636C2DD2A4E3C2D6187E67711F3C8006AD209B5B2161785F36072C92E6E7C24BBB513248AAE60FA240CEBA4E0D96BE865175E262FC97ED063C984C1F8DA1A3264D672F5F62E92BF86319EF59335BF353D6381871BD45C730C2B96CAAC653B01D62C1D9E0261334812A90127648547341F6F740CD14E2CD50606B9CDA91AB", 
x"95DC6F3C2DF2A4E3CBD638EE47715D1C8006AD21195F21417F533632AC92E6E7C24AB75130482BEE0F2241C4BF4E4596BE875165E223BC95E90424D45C17DDA1A3065D853F4F26E98BF80309AF59735973D1963918F17D45C730C2B82CAACE33B01C62C1D9E1261319812F90036EC8747100F6E7C8CD14A28578627BD4DA15C3", 
x"C54C672CA5F2A4E24BD6386E47615F3C8016AD20BB5B21617B573626AC9226C7C24CB3503248ABEE0F2241ACBB0E4D963E075165E262F497ED043C984C1F1DA2A3024DC73F4F2EE90BFC4301AF5973597355963818F13D47C730C2B86CA2C713B014E2C1BDE1261B1001AA900366C8747380B6F740CD14E2CD7C666BDCDA91A7", 
x"C54C6B2EA5D224E2CBD6386CC7715D1C8006AD211B5F204179577632AC92E6E7C24EFF503048ABEE4F2240E4AB4EC5963E86117DEA63F497ED0434944C1789A1A3064DE567573FE92BF8431BEF59735BE341963818713D45C730C3BC6CA04653B0146261DDE126173501AA90127EC85473C0F6F750CD14AACD78622294DA15A3", 
x"97CE6F2D2D92A4E3CBD6386C07715D3C8002AD21395F31615B5F76176C92A6C7C24EFF1032482BE60F2220E4BB0E0D863E86596DE02AF495ED060CC0DC1F9DA1AB035DA73B5F66E98FF40301AF4D735973D1963919F13D47C53082F86C8ACE17B01CE2C19DE1261B1D832F900366C8547140F6E7E8CD14AA8574664A9CDA15A3", 
x"D75C6F2DADF2A4E34BD6387C65715D3C8006AD201B5F31617B5736332C92E6E7C34BFF113248ABEE1FA241C4BF4E4D96BE87196DE262F497ED043CC45C179DA1AB065DE5375723E90BFC6301AF59735973D5D63818713D45C730C3B86C80CE13B09C6241D9E1261B1981AF901376C85471C0B6E740CD14A28558626A9CDA91EB", 
x"855C6F6E2DF2A4E2CBD628EC27715D2C8016AD603B5F376178577632AC92E6C7D34EBB553248ABEE1F2200D4BF4E4586BE87116DE2617C95E9062C845C57DDA4AB075DC537772EE90BFC0301EF5D635973D5D63819713C65C130C2B82CAACF37B0146241D9E1261B15812F80137648FC7340B677E0CD14A29D7C661294DA95E7", 
x"D5CC4B2CADD2A4E3CAF618EC07715D3C8006AD209B5F31617F5F36062C92A6E7C24CF7513248ABEE1FA240C6BF0E4D863E865965E260F495E9063CCC5C575DA1A3264DC52B5F22E9EBFC2301AF5D735BF3D5963818F13D47D73082B92CAACE77B01C62C19DE0261B15812F90027EC85471D2F6F7C0CD14E2857C7262DCDA95A3", 
x"D55C6F6C2DF2A4E3CBD6287C45715D2C8002AD61FB5F374179173632AC12E6E7C34EFB703248ABEE0F2241F4BF4E4D96BE861165C26BF4B5E90438D45C1BCDA2AB074DC5375766E9CBF80303EF4D635D7355D6381971BD65D538C3B964AACF17B09462C1F9E1261B15832E800376C85C7340B267E0CD14A28D5066739CDA95E3", 
x"955C7F2C2DD224E3CBD6287C45715D2C8026AD205B5F346179577632AC92E6C7C34EFF153248ABEE4F2261A6AF4E8D963E871575E262FC97ED0604D05C1B5DA2AB074DC537576EE90BF84301AB4D635F73D5D63019F13D47C730C3B964A84F53B014E2C1D9E1261B1D012F90137648547340B66760DD94A28D5C62739CDA95E3", 
x"C5CC6F6CA5B2A4E28AD6386C47714D3C8006BD21BB5F21617B5736326C92A6E7D24EF7513048ABEE1F2241E6AF460D96BE87136DD022F497E904349C4C17D9A0A30649C72F772FE92BF86309EF49735B7353D63818713D4FC730C3B12CA8CF17B01CE2C19DE0261B3581AE800376C8747380F6E7D8CD14EAC55C7463DCDA95AB", 
x"B54E6F3CADF224E3CAD6187C27715D3C8006BD20795B3061791776076C92E6E7C278FF103248ABE61F2240AEAB468D962E86516DEA68F497AD060C90DC1F1DA0AB024DC5374F73E9EBF46311AF5D735963D5D63919F13C45C73082BD2CAACE57B01D6261FDE1261B3001AE801376C8D471C0F6F7E85D14E2CD7C64629CDA11E3", 
x"954C7F6C2DF2A4E3C3F628FE45715D2C8402AD203B5B356179573637AC9266C7D24FBF513048ABEE4F22C0E4AF0E5D963E86116DC060B497ED063CDCDC57DDA1AB234D25374676E90BFC431BAF5973597355963818717D4FC730C2B86C82CE71B01CEAC1CDE1261B1105AE90036EC8D471C0B66768CD14A2855C62139CDA15E3", 
x"854C6B2EADF2A4E34BD618FE85715D2C8406AD601B5F364179573637AC9266E7D34FBB1032482BE65F22C1C4BF0EDD863E86116FE26AB497A9023AD45C171DA3AB074D8537573EE96BF84303AB5D735F7341D63019715C4FC53082BC64AACE43B01DEAC1DDE1261B15812E90036E48D47340B66760CD14E28D58621B94DA15E3", 
x"87CE4B2CA5F224E34BD638EC25715D3C8002AD21195F3161795736372C92E6C7C24BF75132482BEE5E2240C4BF4E4D863E861165E262B497E9062CDC5C179DA1AB0649A53B5F76E90BD06303EF4D635F73D596B108713C47C730C3B82CA24E11B09DE24199E1261B1901AF901776C85C7340B6E7C0CD14EA8D786262DCDA1583", 
x"F74C7B2C2DF2A4E3CBD638FC45615FAC8006AD603B5F01417C533622EC92E6E7C34BBB713248ABE64E2241B4BF4E0D963E861167E263F495ED0434C85C175DA2A3075DE73F5E67E92BF80309EF49735DF3D1963919F13D45C53883B864A84F17B01CE2C19DE126131181AE90067E485473C0F6F760DD14E2857C627BDCDA15A3", 
x"D9CE6F2C25D2A4E2CBD6186C07715D3C9026BD201B5F34617E5776162C92A6C7C268FB503248ABEE1F2240A4AA460D96AE86596DF261F495ED042CD05C1B0DA1A3024DC52F5F27F9EBF86301AF59335F63C1963919713C45C33082BC6C88CF13B01E6A419DE126131D812E801666C8F473C1F6E760DD14A2CD7C644B9CDA95A3", 
x"D5CC6F6C2DD2A4E34BD6186C47715D3C8016AD203B5B14617D5736262C922647C24AF7503048ABEE4F2241E4BE46CD96BE865165E2697497ED063C944C179DA2A30249C52F5F3EF98BF06301AF5D735963D1963809713D45C738C2B92C80C713B01D62C1BDE1261B1401AE80136EC85C7100B6F760DD14EA8D78647BDCDA91AF", 
x"C74C6F3C2DD224E2CBD6187E6F715F3C9026AD203B5F23617B573636AC92E6E7C359B3503248ABE61F2241E6BA4E0D96BE865365E069F497ED043E984C170DA2A3024DE5275F2BE9EBFC230BAF5963D97353D43108713D45C138C2B964A2CF57B0B4E241FDE1261738092E840276487C73C0F6E7D0CD14A2CD506622DCDA118B", 
x"95DE6B7CADB2A4E3CBD6386C67715D3C8006AD209B5F25617D577612EC12A6E7C25BF3513248ABE60FA240ECBE4E4D96BE861165E263F495ED063CD05C1F0DA1AB0749E52F5F76F9EBFC0303EF59735B73D5963819713C45C338C2B82CA8CE13B03CE241D9E1261B1581AF901376C87C7140B6F740CD14A29D50626BDCDA15E3", 
x"D55E6F2C259224E3CBD6286C67715D9C8002AD60FB5F37417B5736322C1226C7C24AF3513248ABEE0F2241A4BF4ECD86BE871165E268FC97ED0628805C575DA0AB074D85274F36E98FF00311AF5D735D73D5D63009713C45C730C2B96CA84E05B09462C1D9E1261B1101AA801376405C7342B667F0CD14A28D54623394DA1583", 
x"89CC4B6CADB2A4E3CBD6386C47715D3C8002AD203B5F01417F1736062C9226E7C24AFB513248ABEE1F2201ECBF064D96BE875175E269F497ED0628D05C1F19A1A30749E7375F3AF90BF46309AF5D6359F3D1D63919F13D47C73082FD6CA04E33B01C62E199E1261315012A90137EC8D47140F6E770DD14E2CD746479DCDA15AB", 
x"C14C6B6CAD9224E2CAD6386E67715F3C8026AD201B5F34415B5F36226C92E6E7D34AB77130482BEE1F2240ECBB4E0D96BE86577DC26BFC97ED0438984C1F0DA5A3074DE5635726E9ABFC630BAF5D735BF351943919713D47C730C2B96CA24753B03C62E1D9E0261F3481AA80067EC8547381F6E7C0CD14E2CD7C646ADCDA11CB", 
x"915C6F6C2DB2A4E3CAD6287C65715D3C9026AD21B95F31617D5776222C9266E7D24ABF513248AAE60FA200E4BF0E4D86BE861565E222F497E9040CD45C179DA0AB2749A7375E3EE96BFC0301AF4D635B73D5D63919713C47C530C2B924A84753B09C624199E0261B14812F901376C85473C0F6E7F0CD14E2CD7866689CDA95AB", 
x"C15C4B3CADD224E34AD618EC25715D3C8006AD20195B3161795776122C1266C7D25AB7513248ABEE5E2201A4BF0E8D96BE861175EA2BFC95A9063490DC139DA2AB0749853F4F6EF98BF82303AF5D635F73D5D4B918713C67D73882B92CAACE17B03D6A4199E0261B1581AF901766C8FC7102B677705D14E28D54627B9CDA95E3", 
x"E5CC473CADF2A4E24BF6386C67715F3C9036AD603B5B34617D573626AC922647C258B3503248ABEE1FA221A6BE464D96BE865165E0617C97AD0638984C1B1DA5A32749252F5F77E9CBFC6311AF597359F355963109F13C47C13883B96C88C613B01DE2C1DDE1261B3481AE901666C87C7381F6E750DD14E28D706072DCDA91AB", 
x"855E4B2C25F224E3CBD6286C05F15D2C8026AD20DB5F3141795776336C12E6CFD24FFF5132482BEE0F2240A4BF0ECD862E861165C221B495A9062CD45C175DA0AB274DA53B577FE90BF80303EF5D635B73D5963809713C45C738C2FD24A8CE13B03EEAC1D9E1261B1901AF90137E48DC7342B667E0CD14A295587233D4DA15C3", 
x"954C4F2C2DF224E34BD638EC65715D3C9012AD219B5F3161595776132C92A6E7D25EFF513248ABEE4F224184BF4E8586BE87516DE262FCB7ED062CD45C1FDDA0AB0759E53F5767E90BFC6303EB59735963D596B918717D45C738C2B82CA24E13B0966AC1C9E126131581AB90137EC8DC7340B6E748DD14A28D586263D4DA15C3", 
x"954C6B2CADD224E2CBD6386C07714D3C8016AD203B5B20617D5776162C9226C7C34AB7513248ABEE0F2241A4BF46CD96BE86516DE2297C95AD0638944C531DA1A30349E72F5F2EF9CBF84319AB493359E3D1963908713C45C130C3B96C88C633B01D62C1BDE126131089AE80136EC8DC7140F6E760DD14EA8D787673DCDA91E3", 
x"85CE6F2CA5F2A4E34AD6386E05715D3C8006AD60DB5F31417F577626EC92A6E7D24BFF5030482AEE0F2221E4BA064596BE861165E023F497E90638D4DC5719A1A3074DE737562BE9AFF02309EF5D635F73D1D63818F17D4DC73882B96C82C637B01D6AE199E026131D012E900366C8547140F6E7E0DD14AA85786043DCDA95C3", 
x"B5CE6F2F2DD224E3CBD6386E27715D1C8002AD215B5F2441791F36366C9266E7D25BF77132482AEE4F2241CCAF4ECD963E861175E062F4B7ED0634D45C575DA1AB074DE53F7626F92BF8430BAF59735D73D5943818791D45C53083BC2CAACE01B01CE2C1D9E1261F1501AF901376C8547142B6F760DD14A28D5872529CDA15C3", 
x"C5CC4F2C2DF2A4E34BF6186E07715D3C9016BD603B5F35617B5F3607EC92A6E7C248BF5130482BEE0F2241ACBA4E0D96BE06517DF260FC97ED063CD84C1F1DA3A3064DC5275F76E9CBFC2309AB4D735973D1963818F93D47D530C3B86CA84777B01562C19DE1261B3C812E80026EC85C7101B6E7C8DD14A28D70625BDCDA91EB", 
x"C75C6B2E2DD2A4E3CBD6186E27715D3C9006AD215B5F344179137622AC92E6E7C25FBB503248ABE64F2241ACBF4E0D963E86557DE063F497AD0434D85C579DA2AB074DC7277766E9AFD84301AF5D735F63C196B919F13D47D538C3B824A84F03B09CE26199E1261B1081AE900376485C7340B6E760CD14A28D5C664BDCDA95E7", 
x"F14C6F2C2DB2A4E24AD6087E47715D3C8022AD20395F24615D5736066C92E6E7D24EFF513248AAEE1FA260A4AF0E4D86BE86116DD22AF497AD042CD8DC1F5DA0A32749A7275F62E98FFC6319AF49235973D596B918F1BD65C33082B92480CF13B01CE2C199E026133C012E801376C87473C2F6F760CD14A28D74604B9CDA91A3", 
x"854E6F7DADD2A4E34BD6287E67615D3C8022BD21595F00417C573633EC1A62C7C34FB75032482BEE4F2211E4AF4E4D96BE875B75E268F497ED0624D85C1749A1A3074D45377F37F92BDC4303EB5D635D6357D63808713D47D538C3B96CA24E03B0146AE199E1261F1D81AB900376C0547383B66750CD14E2CD7C64439CDA15E3", 
x"C5CC4F2E2DF224E3CBD6386C07F15D3C8026AD20D95F15417B173622EC9266E7C24EFB513248AAEE1F22418CBB4645963E861175EA6BF495E9040C985C171DA3AB0649C7375F2AE92BFC6309AF49635D63D5D4B918F13D45C73082B86CAAC613B01C6AE1D9E1261311012A801366C8FC7340B6F748CD14E28D54624ADCDA15E3", 
x"95CC637CADF2A4E2CAD6186E67714F3C9024BD60BB5F36617D1F36266C92A6C7C358B7503248ABE60F2251E6BB4E45963E875175D063F497ED043E984C1F5DA1AB064DE7235F2AE90BD46303EF5D23596352943018F13D45C338C2B96CA24F17B03DE2C1D9E0261310012E800376C87471C0F6E7D0CD14E2CD78646B9CDA9183", 
x"F54C472CA5B2A4E3CBD6187E47715D3C9026AD20195F11615B577617EC92A6C7C26EF3503248ABE60F2241FCBB460D96BE86116DE262F497ED042CC85C1B1DA1A3075DE73B5F62E9ABF46309AF5D735973D5963919713D65D33082B96CAACE11B01F6261DDE1261318812E90126EC8547341B6E7C8CD14E2C578666B9CDA11A3", 
x"C74C6B2C25F224E34BD6387C07714D2C8026AD215B5F3141795776322C9226E7D24BF7113248ABEE4E224184BF0E4D86BE871165C260FC97AD060CD45C175DA4AB234DC5374F77E96FF00303AD59635F73D196B019F11C47C53082F96CA2C733B01EE2C1D9E1261B19012E90137EC8D47342B66740DD14A2D55C627A94DA1583", 
x"854C7F2C2DF2A4E3CBD6386E07715D2C9006BD61BB5F30417D5F3637AC92E6C7C24BFF5132482AE64F2240A4BB4E4D963E86116DE861F495ED0624C45C135DA1A3274DC53F4F77E92FF86301AF5D735973D5963819F17D47C530C2B96C8A4E51B01CE2C199E1261B1501AE90026EC85473C0F66758CD14E2857076129CDA95E3" 


    );
begin
    process(clk, reset)
    begin
    if (rising_edge(clk)) then
        
        if reset = '1' then
            data_out <= (others => '0'); -- Initialize data_out to zero on reset
        else
            if Read_en = '1' then --when read enable is high
                -- Output 4 bits (one hex digit) from selected address
                -- bit_addr 0 = bits 1023 downto 1020, bit_addr 1 = bits 1019 downto 1016, etc.
                data_out <= ram(to_integer(unsigned(testHV_addr)))((1023 - to_integer(unsigned(bit_addr)) * 4) downto (1020 - to_integer(unsigned(bit_addr)) * 4));
            -- when enable is high, output the corresponding 4-bit hex digit
            --==================
            --When enable is low, do nothing and keep the previous values
            end if;
        end if;
    end if;
    end process;
end Behavioral;