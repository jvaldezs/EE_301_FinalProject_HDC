--------------------------------------------------------------------------------
-- File: ClassHV_RAM.VHD
-- Author: 
-- Date: November 11, 2025
-- Description: RAM module for storing class hypervectors (1024 bits = 256 hex)
--              Sequentially reads out hex values and signals when complete
-- 
-- Revision History:
-- Date          Version     Description
-- 11/11/2025    1.0         Initial creation
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

-- A 1028x26 single-port RAM in VHDL
entity ClassHV_RAM is
port(
 class_select: in std_logic_vector(4 downto 0); -- Select which class (0-25)
 --this input comes from the BIT_SELECT 
 bit_addr: in std_logic_vector(7 downto 0); -- Hex digit address (0-255)
 --this input comes from the BIT_SELECT
 RAM_CLOCK: in std_logic; -- clock input for RAM from top level clock
 RAM_EN: in std_logic; -- Enable reading FROM THE CONTROLLER/STATE MACHINE
 --this input comes from the controller/state machine
 reset: in std_logic; -- Reset input from controller
 RAM_DATA_OUT: out std_logic_vector(1023 downto 0); -- 4-bit hex digit output ** out std_logic_vector(3 downto 0) **
 --data out to the registers feeding the HAMM accumulator
 CLASS_OUT: out std_logic_vector(4 downto 0) -- Output current class being read to the guess compile module

);
end ClassHV_RAM;
architecture Behavioral of ClassHV_RAM is
-- define the new type for the RAM storing hex strings
type RAM_ARRAY is array (0 to 25) of std_logic_vector (1023 downto 0);

-- initial values in the RAM (26 class hypervectors, each 1024 bits)
signal RAM: RAM_ARRAY :=(
x"C54C6F2CADF2A4E3CBD6386C67715D3C8006AD201B5F31617F5736222C92A6E7C24AB7513248ABEE0F2241E4BF4E4D86BE865165E263F497ED063CD05C179DA0AB0749C5375F22E92BF84301AF5D635973D5963819713C45C730C2B92CA8C613B01C624199E1261B1581AE901376C85473C0B6F740CD14A28D58626BDCDA95E3", 
x"D55C6F6CADF224E3CBD6386C05715D2C8006AD201B5F3561795776322C92E6C7D24FBB553248ABEE0F2241E4BF4E4D86BE861165E263F497E90638D45C175DA0AB074DC5375736E9ABF80303AF5D635D73D5D63819713D45C730C3B924A84E13B01CE2C1D9E1261B11012F901366C85C7340B67760CD14A28D58623B9CDA95E3", 
x"85CC6F2C2DD224E3CBD6286E45715D2C8002AD60BB5F35617B573637EC1266C7C34FFF5132482BE60F2240E4AF4ECD863E87116DE062F497ED063CC45C175DA1AB274D85375677E92FF84301EB5D735D73D5963818717D47C538C2B86CAACE13B01CE2C1DDE1261B1501AF901366C85C73C2B66740CD14E28D58621B94DA15E3", 
x"D55C6F6EADD224E3CBD6286C25715D3C8002AD201B5F3561795736322C9266C7D34FFF553248ABEE0F2240C4BF4E4D86BE861165E263F497E9063CD45C175DA0AB074DC5375736E90BF80303EF5D635D73D5D63819713D45C730C2B96CA84E13B01CE2C1D9E1261B1581AF901366C85C7340B66760CD14A28D58721B94DA15E3", 
x"D55C6F6CADF224E3CBD6286C25715D2C8002AD201B5F3761795776322C9266C7D34FBB553248ABEE0F2240C4BF0E4D86BE871565E263F497E9062CD45C17DDA0AB074DC537573EE92BF80303AF5D635D73D5D63819713D45C530C3B964AA4F17B01CE2C1D9E1261B1581AF901366485C7340B67760CD14A28D58621B94DA95E3", 
x"D5CC6F2CADF2A4E2CBD6186C67715D3C8026BD203B5F01617F5736062C92A6E7C24ABF513248ABE61F2241A4BA464D96BE86116DE261F495AD063CD05C1F1DA1A30649C53F5F22E90BFC6309AF5D7359E3D5963918713D47C33082B86CAACF53B01D62619DE126131D812E901776C87471C0F6F760CD14A28D7C647BDCDA11A3", 
x"D55C6F6CADF2A4E3CBD6286C05715D2C8002AD209B5F3141795776322C92E6C7D34FFF513248ABEE0F2240C4BF4E4D863E871165E262F497E9062CD45C175DA0AB274DE5375676E92BF84303EF5D635D73D5963018F13D45C730C2B82CAACE13B01CE2C1D9E1261B1101AF901376C8547340B66760CD14A28D78721B94DA15A3", 
x"D15C6F2CADF224E3CBD6186C65715D3C8022AD201B5F31617D5736062C92E6E7D24AFF513248ABE60F2240C4BF0E4D86BE861165E262F495A9043CD45C1F5DA0AB064DC53F4F66E98BFC2301AF5D735F73D5D63819713C45C33082B92CAACE13B01C624199E1261B15812E901366C8747340B6F760CD14A28D5C627B9CDA95E3", 
x"C5CC6B2CADF2A4E2CBD6386C67715D3C8016AD203B5F21617F5736262C92A6C7C24AB7503048ABEE0F2241A6BE464D96BE865165E269F497ED063C984C171DA1A30249C5275F2AE90BFC2309AF4D3359F3D1963819713C45C730C3B96CA8C733B01D62C19DE1261B1481AA801376C8547180F6E7C0DD14A28D78646BDCDA91A3", 
x"85CC6F2CADF2A4E3CBD6386C67715D3C8002AD201B5F31617F5736362C92A6E7C24AFF503248ABEE0F2241C4BF4E4D863E865165E263FC95ED062CD05C1F5DA1AB075D853F5F66E92BF84301AF59735973D5963818F13D45C730C2B86CAACE13B01CE2C1DDE1261B1501AE90137EC8547340B6E740CD14A28578724BDCDA15A3", 
x"85CC6F2CADF2A4E3CAD6387C67715D3C8002AD201B5F31617F5736362C92A6E7C24AF7513248ABEE0F2241E4BF4E4D96BE861165E263F497ED063CD85C175DA1AB074DC53F5F66E92BF84301AF5D735973D5963818F13D47C730C2B86CAAC613B01C6241DDE1261B1501AE901376C8547140B6E740CD14A28D78626BDCDA15A3", 
x"C54C6F6CADD2A4E3CBD6386C67715D3C8026AD201B5F2061795736222C92A6E7C24ABB503248ABEE0FA240E4BF4E4D96BE865175E26BF497ED043C904C170DA1A3064DE72B5F26E92BF8630BAF597359E3D1963818713D47C730C2B96CA8CF53B01C62C1D9E126133501AA90127EC85471C0F6E760CD14AACD78646B9CDA91A3", 
x"C5CC6F2C25F2A4E3CAD6386C47715D3C8026AD201B5F21417F5736262C92A6E7C24ABF513248ABEE1F2241E4BF0E4D96BE861165E269F497ED063CD05C171DA1A30749C7275F22E92BF8630BAF59635973D1963819713D45C73082B96CA0C753B01C62E199E1261B35012E901376C85471C0F6E760CD14A28D78644BDCDA15E3", 
x"85CC6F2CADF2A4E3CAD6386C47715D3C8026AD201B5F21617F5736262C92A6E7C24AFF503248ABEE1F2241E4BF4E4D96BE861165E263F497E9063CD85C171DA1A30749C7375F26E92BF82309AF5D635973D5943919713D45C73082B96CAAC613B01C626199E1261B3501AE901376C8547140F6E760CD14A28D7C604BDCDA15E3", 
x"C55C6B7C2DD2A4E2CBD6386C67715D3C8026AD201B5F25617B573632AC92A6E7C25BF3503048ABEE1FA241E4BF4E4D96BE865175E263F497ED063C984C170DA1A3074DE5275726E92BF8630BAF59735BF351963818713D47C730C3B96CAAC713B01462C1D9E1261F1481AA901276C8547380F6F7C0CD14E28D58606B9CDA91EB", 
x"D55C6F2CADF224E3CBD6286C25715D3C8002AD201B5F3161795776322C92E6C7C24FBF513248ABEE0F2240C4BF0E4D86BE861165E263F497E9063CD05C175DA0AB074DC5375F76E92BF80303EF59635D73D5963819713D45C730C2B92CAACE13B01CE2C1D9E1261B11012F901376C85C7340B66760CD14A28D58627B94DA15E3", 
x"85CC6F2E2DF224E3CAD6386E67715D3C8006AD611B5F3041791F36336C92E6E7D34BF73032482BEE0F2241C4BF4E0D963E865165E063F497A9063CD05C175DA1AB074DE53F5626E92BF86301AF59735973D5963818717D45C73083B82CA2CE13B01CE2C1D9E1261B1101AA90137EC85471C2B6E760CD14E28578604BD4DA15C3", 
x"C54C6B6C2DD2A4E2CAD6386C47715F3C8026AD203B5F20617F5F3626AC92A6E7C258B7503248ABEE1F2241E4BA4E0D96BE865365E261F497ED063C984C1F0DA1A3064DC52F5F2AE90BFC6303AF5D3359F3D1963818713D47C730C2B96CA0C713B015E2E1D9E1261B3401AA80127EC87473C0F6E7C0CD14E28D786443DCDA91AB", 
x"95CC6F2CADF2A4E3CBD6186C67715F3C8026BD203B5F21617F5736062C92A6E7C25ABF113248ABE61F2241A4BA460D963E86116DE268B497AD063CD05C1F0DA0AB0649C52F5F62E92BFC6309AF5D735B63D5963919713D45C33082B82CA8CF33B01D62619DE126131D812E901376C85471C0B6E7E0CD14A28D7C646BDCDA11A3", 
x"D55C6F2CADF224E3CBD6286C05715D2C8002AD201B5F3161795736332C9266C7D34FFF513248ABEE0F2240C4BF4E4D86BE871165E263F497E90638C05C175DA0AB274D85375E76E98BF80303EF5D635D73D5963018713D47C730C2B92CAACE13B01CE2C1D9E1261B1101AF901366C85C7340B66760CD14A28558723B94DA15E3", 
x"C55C6F2E2DD224E3CBD6386C67715D3C8002AD201B5F214179173632EC92E6E7D24FFF703248ABEE0F2241E4BF4E4D963E865575E263F497E9063CD85C1F5DA0AB074DC73F5726E92BF80301AF59635973D5963918F13D45C730C3B824AACE13B01CE2C1D9E1261B1101AA901376C85473C0F6F7E0CD14A28D5C604BDCDA15E3", 
x"D55C6F2CADD224E3CBD6387C05715D2C8006AD201B5F3541795776322C92E6C7C24EFF513248ABEE0F2240C4BF4E4D86BE861165E263F497E9063CD45C1F5DA0AB074DC5375776E90BF84301AF5D635D73D5D63819713D45C530C2B824AA4E13B01CE2C1D9E1261B11812F901366C85C7340B67760CD14A28D58623B94DA95E3", 
x"D54C6F6C2DD224E3CBD6386C47715D3C8006AD203B5F21417B573632AC92A6E7C24AF7503248ABEE1F2241E4BF4E0D96BE861165E263F497ED063CD84C171DA1A3074DC5375F36E92BFC430BEF59735973D5963818713D45C73083B96CA8C633B01C62E1DDE1261B1501AE901376C85473C0F6E740CD14A28D78666BDCDA15A3", 
x"91CC6F2CA5D2A4E3CBD6187C67715D3C9026BD201B5F20617F5736062C92E6E7C24AFF503248ABE61F2240A4BA464D96BE86116DE269F495AD043CD05C1F5DA1A3064DC73F5F6AE9ABF46301AF5D735B63D1963919713D45C33082B96CA8CF73B01D62419DE1261315812E901776C87471C0B6E760CD14A28D7C667BDCDA95A3", 
x"D54C6F2CADD2A4E2CBD6186C67615F3C8022AD203B5F31617B573636AC92E6C7C25CB7503248ABE60F2241A6BF4E4D96BE865365E263F497ED043C984C1F1DA3AB024DC7275F7BE90BFC2301AF5973597351943818F13D45C530C2B86CA8CF57B015E2C1DDE1261314812A900376C87C73C0F6F7C0CD14A28D5C666BDCDA91A3", 
x"C5CC6F6CADD224E34BD6386EC5715D2C8002AD60BB5F3561795736336C9266C7C34FFF1132482BEE0F2241E4BF4E4D863E871165E062F497E9063CC45C1F5DA0AB274D85375677E92FF80301EB5D735D73D5D63818713D47C538C2B86CA8CE07B01CE2C1D9E1261B1501AF901366485C73C0B66760CD14E28D58621B94DA95E3" 


   ); 
begin 
    process(RAM_CLOCK, reset)
    begin
    if(rising_edge(RAM_CLOCK)) then
        if(reset = '1') then
        -- Reset the RAM data output 
        
            RAM_DATA_OUT <= (others => '1'); -- Initialize data_out to zero on reset
        elsif(RAM_EN = '1') then --should be controlled by controller/state
        -- Output 4 bits (one hex digit) from selected class at specified hex digit address
        -- bit_addr 0 = bits 1023 downto 1020, bit_addr 1 = bits 1019 downto 1016, etc.
        RAM_DATA_OUT <= RAM(to_integer(unsigned(class_select)));
        --address is selected by the class and the bit_addr input and uses the above function to call the individual binary bits of each individual hex bit since the array is indexed as...
        -- hex making the individual bits avialable to access from 0-1023
        -- RAM_DATA_OUT <= RAM(to_integer(unsigned(class_select)))((1023 - to_integer(unsigned(bit_addr)) * 4) downto (1020 - to_integer(unsigned(bit_addr)) * 4));
        end if;
        -- Always output the current class select (combinational, not gated by RAM_EN)
        CLASS_OUT <= class_select;
    end if;
end process;

end Behavioral; 

